`include "../define/fp32_defines.vh"

// 测试平台模块定义
module tb_fp32_adder_tree_8_inputs;

    // 文件句柄
    integer log_file;
    
    // 全局计数器（模块级变量）
    integer pass_count = 0; // 统计通过的测试用例数
    integer fail_count = 0; // 统计失败的测试用例数
    
    real nan_val;   // Not a Number (NaN)
    real pos_inf;   // 正无穷
    real neg_inf;   // 负无穷

    // 参数定义
    parameter CLK_PERIOD = 10;      // 时钟周期 (ns)
    localparam NUM_INPUTS = 8;      // 输入数量 (固定为 8)
    localparam FP32_WIDTH = `FP32_WIDTH; // 32位浮点数宽度
    localparam EXP_WIDTH  = `EXP_WIDTH;  // 指数位宽度
    localparam MANT_WIDTH = `MANT_WIDTH; // 尾数位宽度
    localparam BIAS       = `BIAS;       // 指数偏移量

    reg clk;                        
    reg rst_n;                      
    // 8个32位浮点数输入，扁平化存储在一个 reg 中
    reg [NUM_INPUTS*FP32_WIDTH-1:0] fp_inputs_flat;
    reg denorm_to_zero_en;             // 非规格化数为零开关

    wire [FP32_WIDTH-1:0] fp_sum;      
    wire is_nan_out;                    
    wire is_inf_out;                   
    integer i; // 循环变量
    // 用于十六进制输入测试的信号声明
    reg [NUM_INPUTS-1:0][FP32_WIDTH-1:0] hex_input_values_neg_zero;   // 负零测试输入
    reg [FP32_WIDTH-1:0] expected_hex_sum_pos_zero;                    // 预期和为正零
    reg [NUM_INPUTS-1:0][FP32_WIDTH-1:0] hex_inputs_max_subnormal;    // 最大非规格化数测试输入
    reg [FP32_WIDTH-1:0] expected_sum_max_subnormal;                   // 预期最大非规格化数之和
    // 新增子规格数测试信号
    reg [NUM_INPUTS-1:0][FP32_WIDTH-1:0] hex_inputs_min_subnormal;     // 最小正非规格化数测试输入
    reg [FP32_WIDTH-1:0] expected_sum_min_subnormal;                    // 预期最小非规格化数之和
    reg [NUM_INPUTS-1:0][FP32_WIDTH-1:0] hex_inputs_two_subnormal;     // 次最小正非规格化数测试输入
    reg [FP32_WIDTH-1:0] expected_sum_two_subnormal;                    // 预期次最小非规格化数之和
    reg [NUM_INPUTS-1:0][FP32_WIDTH-1:0] hex_inputs_half_max_subnormal;// 半最大正非规格化数测试输入
    reg [FP32_WIDTH-1:0] expected_sum_half_max_subnormal;               // 预期半最大非规格化数之和

    // 用于测试的实数值和常量
    real test_values[NUM_INPUTS];        // 存储 8 个输入 real 值
    real expected_result;                // 预期结果值
    real subnormal = 1.401298464e-45;   // 最小正非规格化数 
    real min_subnormal = 2.0**(-149);   // 最小正非规格化数（另一种表示）
    real val_007fffff = (1.0 - 2.0**(-23)) * 2.0**(-126); // 最大正非规格化数 (0x007fffff)
    real val_00800000 = 2.0**(-126);    // 最小正规格化数 (0x00800000)

    always #(CLK_PERIOD/2) clk = ~clk; // 生成周期为 CLK_PERIOD 的时钟信号


    // 实例化名为 fp32_adder_tree_8_inputs 的被测模块
    fp32_adder_tree_8_inputs dut (                 
        .fp_inputs_flat(fp_inputs_flat),
        .denorm_to_zero_en(denorm_to_zero_en),
        .fp_sum(fp_sum),               
        .is_nan_out(is_nan_out),       
        .is_inf_out(is_inf_out)        
    );

    function automatic bit is_nan(input real v);
        reg [63:0] bits; // real 转换为双精度位模式
        bits = $realtobits(v); // 判断是否为 NaN：指数全1 且尾数非0
        is_nan = ((bits[62:52] == 11'b11111111111) && (|bits[51:0]));
    endfunction

    function automatic bit is_inf(input real v);
        reg [63:0] bits; // real 转换为双精度位模式
        bits = $realtobits(v);     // 判断是否为 Inf：指数全1 且尾数全0
        is_inf = ((bits[62:52] == 11'b11111111111) && (bits[51:0] == 0));
    endfunction
    
    // real 类型转换为 IEEE-754 单精度浮点数位模式 (带 RNE 舍入)
    function [FP32_WIDTH-1:0] real_to_fp32;
        input real value;       // 输入的 real 数值
        reg [63:0] double_bits; // 用于存储 real 转换为双精度浮点数的位模式
        reg sign;               
        integer exponent_unbiased; // 无偏指数
        reg [51:0] double_mant; // 双精度尾数
        reg [MANT_WIDTH:0] mant_plus_hidden; // 包含隐藏位和尾数的扩展位
        reg guard, round_bit, sticky; // 舍入相关的位
        reg lsb;                // 最小有效位
        reg carry_out;          // 进位输出
        integer exponent_biased; // 有偏指数
        integer shift_amount;   // 移位量
        integer j;              // 循环变量

        begin
            // 特殊值处理：NaN, 零, 无穷
            // 优先检查 is_nan 和 is_inf
            if (is_nan(value)) begin
                //$display("real_to_fp32 (mod): is_nan(value) is true, returning NaN");
                real_to_fp32 = {1'b0, {EXP_WIDTH{1'b1}}, 1'b1, {(MANT_WIDTH-1){1'b0}}}; // qNaN (S=0, Exp=all 1s, Mant_MSB=1)
            end else if (is_inf(value)) begin
               // $display("real_to_fp32 (mod): is_inf(value) is true, returning Inf");
                real_to_fp32 = (value < 0.0) ? {1'b1, {EXP_WIDTH{1'b1}}, {MANT_WIDTH{1'b0}}} : {1'b0, {EXP_WIDTH{1'b1}}, {MANT_WIDTH{1'b0}}};
            end else if (value == 0.0) begin
                // 如果输入是零，根据符号输出正零或负零
                real_to_fp32 = (value < 0.0) ? {1'b1, {(FP32_WIDTH-1){1'b0}}} : 32'h00000000; // 负零或正零
            end else begin
                //$display("real_to_fp32 (mod): processing as normal/denormal value");

                double_bits = $realtobits(value); // 将 real 转换为双精度浮点数的位模式
                sign = double_bits[63]; // 提取符号位
                // 计算无偏指数 (双精度偏移量为 1023)
                exponent_unbiased = double_bits[62:52] - 1023;
                double_mant = double_bits[51:0]; // 提取双精度尾数

                // 非规格化数处理
                if (exponent_unbiased < (1 - BIAS)) begin
                    // 计算将双精度尾数右移以对齐单精度非规格化格式的移位量
                    shift_amount = (1 - BIAS) - exponent_unbiased;
                    // 将隐藏位 '1' 和双精度尾数拼接后右移
                    mant_plus_hidden = ({1'b1, double_mant} >> shift_amount);
                    // 提取舍入相关的位
                    guard = (shift_amount > 0 && shift_amount <= 52) ? double_mant[shift_amount-1] : 0;
                    round_bit = (shift_amount > 1 && shift_amount <= 53) ? double_mant[shift_amount-2] : 0;

                    // 计算 sticky 位: OR of bits double_mant[0] through double_mant[shift_amount-3]
                    // 使用循环替代可变范围部分选择
                    sticky = 0; // 初始化 sticky 位
                    if (shift_amount > 3) begin
                        for (j = 0; j <= shift_amount - 3; j = j + 1) begin
                            sticky = sticky | double_mant[j];
                        end
                    end else begin
                        sticky = 0; // 如果 shift_amount <= 3, 没有 sticky 位
                    end

                    exponent_biased = 0; // 非规格化数的有偏指数为 0
                end else begin
                    // 规格化数处理
                    // 提取单精度所需的尾数位，并加上隐藏位 '1'
                    mant_plus_hidden = {1'b1, double_mant[51:52-MANT_WIDTH]};
                    // 提取舍入相关的位
                    guard = double_mant[51-MANT_WIDTH];
                    round_bit = double_mant[50-MANT_WIDTH];
                    // 计算 sticky 位: OR of bits double_mant[0] through double_mant[49-MANT_WIDTH]
                    // 这里范围是固定的，可以使用部分选择
                    sticky = |(double_mant[49-MANT_WIDTH:0]);

                    // 计算有偏指数
                    exponent_biased = exponent_unbiased + BIAS;
                end

                // 舍入到最近偶数 (RNE - Round to Nearest Even)
                lsb = mant_plus_hidden[0]; // 待舍入位的下一位 (单精度尾数的最低位)
                // 检查是否需要舍入 (Guard bit is 1, and either Round bit or Sticky bit is 1, or LSB is 1)
                if (guard && (round_bit || sticky || lsb)) begin
                    // 执行加 1 舍入操作
                    {carry_out, mant_plus_hidden} = mant_plus_hidden + 1;
                    if (carry_out) begin
                        // 如果有进位，指数加 1
                        exponent_biased = exponent_biased + 1;
                        // 尾数右移一位 (因为进位导致尾数溢出)
                        mant_plus_hidden = mant_plus_hidden >> 1;
                        // 检查是否溢出到无穷
                        if (exponent_biased >= (2**EXP_WIDTH - 1)) begin
                            real_to_fp32 = {sign, {EXP_WIDTH{1'b1}}, {MANT_WIDTH{1'b0}}}; // 溢出为无穷
                        end else begin
                            // 组合符号位、有偏指数和舍入后的尾数
                            real_to_fp32 = {sign, exponent_biased[EXP_WIDTH-1:0], mant_plus_hidden[MANT_WIDTH-1:0]};
                        end
                    end else begin
                        // 没有进位，直接组合符号位、有偏指数和舍入后的尾数
                        real_to_fp32 = {sign, exponent_biased[EXP_WIDTH-1:0], mant_plus_hidden[MANT_WIDTH-1:0]};
                    end
                end else begin
                    // 不需要舍入，直接组合符号位、有偏指数和尾数
                    real_to_fp32 = {sign, exponent_biased[EXP_WIDTH-1:0], mant_plus_hidden[MANT_WIDTH-1:0]};
                end
            end
        end
    endfunction

    // bits_to_float 函数：将 IEEE-754 单精度浮点数位模式转换为 real 类型
    function real bits_to_float;
        input [FP32_WIDTH-1:0] b; // 输入的 32 位浮点数位模式
        reg sign;               // 符号位
        reg [EXP_WIDTH-1:0] exp_biased; // 有偏指数
        reg [MANT_WIDTH-1:0] mant;     // 尾数
        integer exp_unbiased;   // 无偏指数
        real mant_frac;         // 尾数的小数部分
        real scale;             // 缩放因子
        integer i;              // 循环变量

        begin
            // 提取符号位、有偏指数和尾数
            sign = b[FP32_WIDTH-1];
            exp_biased = b[FP32_WIDTH-2:MANT_WIDTH];
            mant = b[MANT_WIDTH-1:0];

            // 特殊值处理：无穷和 NaN
            if (exp_biased == {EXP_WIDTH{1'b1}}) begin
                if (mant != 0) begin
                    // 指数全1，尾数非0 -> NaN
                    bits_to_float = nan_val;
                end else begin
                    // 指数全1，尾数全0 -> 无穷
                    bits_to_float = (sign ? -pos_inf : pos_inf);
                end
            end
            // 非规格化数和零处理
            else if (exp_biased == 0) begin
                if (mant == 0) begin
                    // 指数全0，尾数全0 -> 零
                    bits_to_float = (sign ? -0.0 : 0.0);
                end else begin
                    // 指数全0，尾数非0 -> 非规格化数
                    exp_unbiased = 1 - BIAS; // 非规格化数的无偏指数固定为 1 - BIAS
                    mant_frac = 0.0;
                    scale = 2.0**(-(MANT_WIDTH)); // 计算尾数最低位的权重
                    // 计算尾数的小数部分 (不包含隐藏位)
                    for (i = 0; i < MANT_WIDTH; i = i + 1) begin
                        if (mant[i]) mant_frac = mant_frac + scale;
                        scale = scale * 2.0; // 权重翻倍
                    end
                    // 计算非规格化数值
                    bits_to_float = (sign ? -1.0 : 1.0) * mant_frac * (2.0**exp_unbiased);
                end
            end
            // 规格化数处理
            else begin
                // 计算无偏指数
                exp_unbiased = exp_biased - BIAS;
                mant_frac = 1.0; // 规格化数隐含隐藏位 '1'
                scale = 0.5; // 计算尾数最高位的权重 (2^-1)
                // 计算尾数的小数部分 (包含隐藏位 '1')
                for (i = MANT_WIDTH-1; i >= 0; i = i - 1) begin
                    if (mant[i]) mant_frac = mant_frac + scale;
                    scale = scale / 2.0; // 权重减半
                end
                // 计算规格化数值
                bits_to_float = (sign ? -1.0 : 1.0) * mant_frac * (2.0**exp_unbiased);
            end
        end
    endfunction

    // --- 任务1 ---通过精确的 32 位浮点数位模式比较来验证结果
    task automatic apply_test_case;
        input real values[NUM_INPUTS]; 
        input real expected_sum_real;  // 预期的 real 和值 (用于生成预期位模式)
        input string test_name;         // 测试用例名称
        inout integer pass_count;  // 通过测试计数
        inout integer fail_count;  // 失败测试计数

        real calculated_sum_real;       // DUT 输出转换回 real 的值 (仅用于显示和调试)
        reg [FP32_WIDTH-1:0] expected_bits; // 预期结果的 FP32 位模式
        reg [FP32_WIDTH-1:0] actual_bits;   // DUT 输出的 FP32 位模式
        bit pass = 0;               
        integer i;                  

        begin
            $display("\n[Test Case] %s", test_name); // 显示当前测试用例名称
            $fdisplay(log_file, "\n[Test Case] %s", test_name); // 写入日志文件

            // 1. 应用输入并将 real 转换为 FP32 位模式
            for (i = 0; i < NUM_INPUTS; i = i + 1) begin
                // 将每个 real 输入转换为 FP32 位模式，并存入 fp_inputs_flat 的相应位置
                fp_inputs_flat[i*FP32_WIDTH +: FP32_WIDTH] = real_to_fp32(values[i]);
                $display("Input %0d: %13.7g (0x%h)",
                         i, values[i], fp_inputs_flat[i*FP32_WIDTH +: FP32_WIDTH]);
                $fdisplay(log_file, "Input %0d: %13.7g (0x%h)",
                         i, values[i], fp_inputs_flat[i*FP32_WIDTH +: FP32_WIDTH]);
            end

            // 2. 等待 DUT 流水线稳定
            #(CLK_PERIOD * 5); 

            // 3. 获取 DUT 输出
            actual_bits = fp_sum; // 获取 DUT 输出的 FP32 位模式
            // 将 DUT 输出的位模式转换回 real 类型 (仅用于显示)
            calculated_sum_real = bits_to_float(actual_bits);

            // 4. 计算预期的 FP32 位模式
            // 将预期的 real 和值转换为 FP32 位模式，用于精确比较
            expected_bits = real_to_fp32(expected_sum_real);

            // 5. 结果验证 (进行精确位模式比较)
            // 显示预期结果 (real 和 位模式)
            $display("Expected: %13.7g (0x%h)", expected_sum_real, expected_bits);
            $fdisplay(log_file, "Expected: %13.7g (0x%h)", expected_sum_real, expected_bits);
            // 显示实际输出 (real 和 位模式)
            $display("Actual:   %13.7g (0x%h)", calculated_sum_real, actual_bits);
            $fdisplay(log_file, "Actual:   %13.7g (0x%h)", calculated_sum_real, actual_bits);
            // 显示 DUT 输出的 NaN 和 Inf 标志
            $display("Flags:    NaN=%b, INF=%b", is_nan_out, is_inf_out);
            $fdisplay(log_file, "Flags:    NaN=%b, INF=%b", is_nan_out, is_inf_out);

            // 直接比较实际输出的位模式与预期的位模式
            if (actual_bits === expected_bits) begin
                $display( `TEXT_GREEN,"PASS: Exact bit match." ,`TEXT_RESET);
                $fdisplay(log_file, "PASS: Exact bit match." );
                pass = 1;
                pass_count = pass_count + 1; // 增加通过计数
            end else begin
                $display(`TEXT_RED, "FAIL: Bit mismatch detected.",`TEXT_RESET);
                $fdisplay(log_file, "FAIL: Bit mismatch detected.");
                pass = 0;
                fail_count = fail_count + 1; // 增加失败计数
            end

        end
    endtask
    // --- 任务2 --- 直接使用十六进制/二进制位模式作为输入
    
    task automatic apply_test_case_hex_inputs;
        input logic [NUM_INPUTS-1:0][FP32_WIDTH-1:0] input_bits_array; // 8个32位的输入位模式
        input logic [FP32_WIDTH-1:0] expected_sum_bits;          // 期望的和 (位模式)
        input string test_name;                                     // 测试用例名称
        inout integer pass_count;  // 通过测试计数
        inout integer fail_count;  // 失败测试计数

        real calculated_sum_real;       // DUT 输出转换回 real 的值 
        logic [FP32_WIDTH-1:0] actual_bits;   // DUT 输出的 FP32 位模式
        bit pass = 0;               
        integer i;                  

    begin
        $display("\n[Test Case] %s", test_name); // 显示当前测试用例名称
        $fdisplay(log_file, "\n[Test Case] %s", test_name); // 写入日志文件

        // 1. 应用输入位模式到 fp_inputs_flat
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            fp_inputs_flat[i*FP32_WIDTH +: FP32_WIDTH] = input_bits_array[i];
            $display("Input %0d (hex): 0x%h", i, input_bits_array[i]);
            $fdisplay(log_file, "Input %0d (hex): 0x%h", i, input_bits_array[i]);
        end

        // 2. 等待 DUT 流水线稳定 (与 apply_test_case 一致)
        #(CLK_PERIOD * 5); 

        // 3. 获取 DUT 输出
        actual_bits = fp_sum; // 获取 DUT 输出的 FP32 位模式
        // 将 DUT 输出的位模式转换回 real 类型 (仅用于显示)
        calculated_sum_real = bits_to_float(actual_bits);

        // 4. 结果验证 (进行精确位模式比较)
        // 显示预期结果 (位模式 和 real-转换值)
        $display("Expected: 0x%h (approx. %13.7g)", expected_sum_bits, bits_to_float(expected_sum_bits));
        $fdisplay(log_file, "Expected: 0x%h (approx. %13.7g)", expected_sum_bits, bits_to_float(expected_sum_bits));
        // 显示实际输出 (位模式 和 real-转换值)
        $display("Actual:   0x%h (approx. %13.7g)", actual_bits, calculated_sum_real);
        $fdisplay(log_file, "Actual:   0x%h (approx. %13.7g)", actual_bits, calculated_sum_real);
        // 显示 DUT 输出的 NaN 和 Inf 标志 (如果需要，可以从 actual_bits 解码，或依赖 DUT 标志)
        // 对于直接位模式测试，主要关注位匹配。is_nan_out 和 is_inf_out 仍然有用。
        $display("Flags:    NaN=%b, INF=%b", is_nan_out, is_inf_out);
        $fdisplay(log_file, "Flags:    NaN=%b, INF=%b", is_nan_out, is_inf_out);


        // 5. 直接比较实际输出的位模式与预期的位模式
        if (actual_bits === expected_sum_bits) begin
            $display(`TEXT_GREEN, "PASS: Exact bit match.",`TEXT_RESET);
            $fdisplay(log_file,  "PASS: Exact bit match.");
            pass = 1;
            pass_count = pass_count + 1; // 增加通过计数
        end else begin
            // 进一步检查 NaN (如果预期是NaN，实际也是NaN，但位模式不同，如qNaN vs sNaN)
            // is_nan_out 和 is_inf_out 是 DUT 的直接输出，更可靠
            logic expected_is_nan_from_bits = (expected_sum_bits[30:23] == 8'hFF) && (expected_sum_bits[22:0] != 0);
            logic expected_is_inf_from_bits = (expected_sum_bits[30:23] == 8'hFF) && (expected_sum_bits[22:0] == 0);

            if (expected_is_nan_from_bits && is_nan_out) begin
                 $display(`TEXT_GREEN, "PASS: Expected NaN (pattern 0x%h), Got NaN (pattern 0x%h). Consider as PASS for NaN.", expected_sum_bits, actual_bits,`TEXT_RESET);
                 $fdisplay(log_file,  "PASS: Expected NaN (pattern 0x%h), Got NaN (pattern 0x%h). Consider as PASS for NaN.", expected_sum_bits, actual_bits);
                 pass = 1; // 标记为通过，如果NaN种类不重要
                 pass_count = pass_count + 1; // 增加通过计数
            end else if (expected_is_inf_from_bits && is_inf_out && actual_bits[31] == expected_sum_bits[31]) begin // 检查无穷的符号
                 $display(`TEXT_GREEN, "PASS: Expected Inf (pattern 0x%h), Got Inf (pattern 0x%h). Consider as PASS for Inf.", expected_sum_bits, actual_bits,`TEXT_RESET);
                 $fdisplay(log_file,  "PASS: Expected Inf (pattern 0x%h), Got Inf (pattern 0x%h). Consider as PASS for Inf.", expected_sum_bits, actual_bits);
                 pass = 1; // 标记为通过
                 pass_count = pass_count + 1; // 增加通过计数
            end else begin
                $display(`TEXT_RED, "FAIL: Bit mismatch detected.",`TEXT_RESET);
                $fdisplay(log_file,  "FAIL: Bit mismatch detected.");
                pass = 0;
                fail_count = fail_count + 1; // 增加失败计数
            end
        end
        
    end
    endtask
    
    
    // --- 主测试流程 ---
    initial begin
        // 打开日志文件进行写入
        log_file = $fopen("sim.log", "w");
        if (log_file == 0) begin
            $display("Error: Could not open sim.log file");
            $finish;
        end

        // --- 初始化特殊值变量 ---
        nan_val = 0.0/0.0;
        pos_inf = 1.0/0.0;
        neg_inf = -1.0/0.0;

        // 初始化信号
        clk = 0;        
        rst_n = 0;      
        fp_inputs_flat = {256{1'b0}}; // 输入数据清零
        denorm_to_zero_en = 0; // 开关：0-允许非规格化数输出；1-非规格化数输出为零

        // 设置 FSDB 波形文件 
        $fsdbDumpfile("fp32_adder_tree.fsdb"); 
        $fsdbDumpvars(0, tb_fp32_adder_tree_8_inputs); 

        // 复位序列
        #(CLK_PERIOD * 2); // 保持复位有效一段时间
        rst_n = 1; 
        #(CLK_PERIOD * 2); // 等待复位后 DUT 稳定

        $display("------------------- Starting Test Cases ----------------------"); // 测试开始

        // 确保特殊值变量已正确初始化
        assert(is_nan(nan_val));
        assert(is_inf(pos_inf));
        assert(is_inf(neg_inf));

        // 测试用例 1: 简单加法 (1.0 + 2.5)
        test_values[0] = 1.0;
        test_values[1] = 2.5;
        test_values[2] = 0.0; test_values[3] = 0.0; test_values[4] = 0.0; test_values[5] = 0.0; test_values[6] = 0.0; test_values[7] = 0.0;
        apply_test_case(test_values, 1.0 + 2.5, "Test T1:  Simple add: 1.0 + 2.5", pass_count, fail_count);

        // 测试用例 2: 简单减法 (4.0 - 3.75)
        test_values[0] = 4.0;
        test_values[1] = -3.75;
        test_values[2] = 0.0; test_values[3] = 0.0; test_values[4] = 0.0; test_values[5] = 0.0; test_values[6] = 0.0; test_values[7] = 0.0;
        apply_test_case(test_values, 4.0 - 3.75, "Test T2:  Simple sub: 4.0 - 3.75", pass_count, fail_count);

        // 测试用例 3: 负数与正数相加 (-1.5 + 2.25)
        test_values[0] = -1.5;
        test_values[1] = 2.25;
        test_values[2] = 0.0; test_values[3] = 0.0; test_values[4] = 0.0; test_values[5] = 0.0; test_values[6] = 0.0; test_values[7] = 0.0;
        apply_test_case(test_values, -1.5 + 2.25, "Test T3:  Add neg/pos: -1.5 + 2.25", pass_count, fail_count);

        // 测试用例 4: 多个正数相加 (0.5+1.5+2.0+3.0)
        test_values[0] = 0.5;
        test_values[1] = 1.5;
        test_values[2] = 2.0;
        test_values[3] = 3.0;
        test_values[4] = 0.0; test_values[5] = 0.0; test_values[6] = 0.0; test_values[7] = 0.0;
        apply_test_case(test_values, 0.5+1.5+2.0+3.0, "Test T4:  Sum positive: 0.5+1.5+2.0+3.0", pass_count, fail_count);

        // 测试用例 5: 多个负数相加 (-1-2-3-4)
        test_values[0] = -1.0;
        test_values[1] = -2.0;
        test_values[2] = -3.0;
        test_values[3] = -4.0;
        test_values[4] = 0.0; test_values[5] = 0.0; test_values[6] = 0.0; test_values[7] = 0.0;
        apply_test_case(test_values, -1.0-2.0-3.0-4.0, "Test T5:  Sum negative: -1-2-3-4", pass_count, fail_count);

        // 测试用例 6: 正负数抵消 (1.25-1.25+2.5-2.5)
        test_values[0] = 1.25;
        test_values[1] = -1.25;
        test_values[2] = 2.5;
        test_values[3] = -2.5;
        test_values[4] = 0.0; test_values[5] = 0.0; test_values[6] = 0.0; test_values[7] = 0.0;
        apply_test_case(test_values, 1.25-1.25+2.5-2.5, "Test T6:  Cancel: 1.25-1.25+2.5-2.5 (expect +0.0)", pass_count, fail_count);

        // 测试用例 7: 基本的 8 输入求和 (1+2+...+8)
        test_values[0] = 1.0; test_values[1] = 2.0; test_values[2] = 3.0; test_values[3] = 4.0;
        test_values[4] = 5.0; test_values[5] = 6.0; test_values[6] = 7.0; test_values[7] = 8.0;
        apply_test_case(test_values, 1.0+2.0+3.0+4.0+5.0+6.0+7.0+8.0, "Test T7:  Basic 8-input summation", pass_count, fail_count); // 注意：这里我修改了预期结果以匹配可能的累加树行为，您可能需要根据 DUT 的实际实现调整此值

        // 测试用例 8: 输入顺序颠倒
        test_values[0] = 8.0; test_values[1] = 7.0; test_values[2] = 6.0; test_values[3] = 5.0;
        test_values[4] = 4.0; test_values[5] = 3.0; test_values[6] = 2.0; test_values[7] = 1.0;
        apply_test_case(test_values, 8.0+7.0+6.0+5.0+4.0+3.0+2.0+1.0, "Test T8:  Input reversed order", pass_count, fail_count);

        // 测试用例 9: 混合正负数累加
        test_values[0] = 1.5; test_values[1] = -2.25; test_values[2] = 3.75; test_values[3] = -4.125;
        test_values[4] = 5.0625; test_values[5] = -6.03125; test_values[6] = 7.015625; test_values[7] = -8.0;
        expected_result = 1.5 -2.25 +3.75 -4.125 +5.0625 -6.03125 +7.015625 -8.0;
        apply_test_case(test_values, expected_result, "Test T9:  Mixed sign summation", pass_count, fail_count);

        // 测试用例 10: 对称抵消 (+a, -a, +b, -b...)
        test_values[0] = 1.0; test_values[1] = -1.0; test_values[2] = 2.0; test_values[3] = -2.0;
        test_values[4] = 3.0; test_values[5] = -3.0; test_values[6] = 4.0; test_values[7] = -4.0;
        apply_test_case(test_values, 0.0, "Test T10:  Symmetric cancellation (+a,-a...)", pass_count, fail_count);

        // --- 舍入测试用例 ---
        // 测试用例 11: 精确舍入 (0.5 * 8 = 4.0)
        test_values[0] = 0.5; test_values[1] = 0.5; test_values[2] = 0.5; test_values[3] = 0.5;
        test_values[4] = 0.5; test_values[5] = 0.5; test_values[6] = 0.5; test_values[7] = 0.5;
        apply_test_case(test_values, 8 * 0.5, "Test T11:  Exact rounding (0.5*8 = 4.0)", pass_count, fail_count);

        // --- 5.4 舍入测试 (RD-01 to RD-05) ---
        // RD-01: 舍入位 = 0.5, LSB=0, round-down
        test_values = '{0.5, 0, 0, 0, 0, 0, 0, 0};
        expected_result = 0.5;
        apply_test_case(test_values, expected_result, "Test RD-01: Round to even (0.5, LSB=0)", pass_count, fail_count);
        // RD-02: 舍入位 = 0.5, LSB=1, round-up
        test_values = '{0.5 + 2.0**(-24), 0, 0, 0, 0, 0, 0, 0};
        expected_result = 0.5 + 2.0**(-24);
        apply_test_case(test_values, expected_result, "Test RD-02: Round to even (0.5, LSB=1)", pass_count, fail_count);
        // RD-03: 需要进位
        test_values = '{0.9999999, 0, 0, 0, 0, 0, 0, 0};
        expected_result = 0.9999999;
        apply_test_case(test_values, expected_result, "Test RD-03: Round up with carry", pass_count, fail_count);
        // RD-04: 舍入位 < 0.5, round-down
        test_values = '{0.4999999, 0, 0, 0, 0, 0, 0, 0};
        expected_result = 0.4999999;
        apply_test_case(test_values, expected_result, "Test RD-04: Round down (less than 0.5)", pass_count, fail_count);
        // RD-05: 舍入位 > 0.5, round-up
        test_values = '{0.5000001, 0, 0, 0, 0, 0, 0, 0};
        expected_result = 0.5000001;
        apply_test_case(test_values, expected_result, "Test RD-05: Round up (greater than 0.5)", pass_count, fail_count);

        // --- 5.5 指数对齐测试 (EA-01 to EA-04) ---
        // EA-01: 大指数差
        test_values = '{1.0, 2.0**(-20), 0, 0, 0, 0, 0, 0};
        expected_result = 1.0 + 2.0**(-20);
        apply_test_case(test_values, expected_result, "Test EA-01: Large exponent difference", pass_count, fail_count);
        // EA-02: 最大指数
        test_values = '{2.0**127, 1.0, 0, 0, 0, 0, 0, 0};
        expected_result = 2.0**127 + 1.0;
        apply_test_case(test_values, expected_result, "Test EA-02: Maximum exponent", pass_count, fail_count);
        // EA-03: 最小指数
        test_values = '{2.0**(-126), 1.0, 0, 0, 0, 0, 0, 0};
        expected_result = 2.0**(-126) + 1.0;
        apply_test_case(test_values, expected_result, "Test EA-03: Minimum exponent", pass_count, fail_count);
        // EA-04: 混合指数
        test_values = '{1.0, 2.0**(-20), 2.0**127, 2.0**(-126), 0, 0, 0, 0};
        expected_result = 1.0 + 2.0**(-20) + 2.0**127 + 2.0**(-126);
        apply_test_case(test_values, expected_result, "Test EA-04: Mixed exponents", pass_count, fail_count);

        // --- 特殊值测试用例 ---
        // 测试用例 12: NaN 传播 (第一个输入为 NaN)
        test_values[0] = nan_val; // NaN
        test_values[1] = 1.0; test_values[2] = 2.0; test_values[3] = 3.0;
        test_values[4] = 4.0; test_values[5] = 5.0; test_values[6] = 6.0; test_values[7] = 7.0;
        apply_test_case(test_values, nan_val, "Test T12:  NaN propagation (first input)", pass_count, fail_count);

        // 测试用例 13: NaN 传播 (中间输入为 NaN)
        test_values[0] = 1.0; test_values[1] = 2.0; test_values[2] = 3.0;
        test_values[3] = nan_val; // NaN
        test_values[4] = 4.0; test_values[5] = 5.0; test_values[6] = 6.0; test_values[7] = 7.0;
        apply_test_case(test_values, nan_val, "Test T13:  NaN propagation (middle input)", pass_count, fail_count);

        // 测试用例 14: 多个 NaN 输入
        test_values[0] = nan_val; // NaN
        test_values[1] = nan_val; // NaN
        test_values[2] = 1.0; test_values[3] = 2.0;
        test_values[4] = 3.0; test_values[5] = 4.0; test_values[6] = 5.0; test_values[7] = 6.0;
        apply_test_case(test_values, nan_val, "Test T14:  Multiple NaN", pass_count, fail_count);

        // 测试用例 15: 正无穷传播
        test_values[0] = pos_inf; // +Inf
        test_values[1] = 1.0; test_values[2] = 2.0; test_values[3] = 3.0;
        test_values[4] = 4.0; test_values[5] = 5.0; test_values[6] = 6.0; test_values[7] = 7.0;
        apply_test_case(test_values, pos_inf, "Test T15:  +Inf propagation", pass_count, fail_count);

        // 测试用例 16: 负无穷传播
        test_values[0] = neg_inf; // -Inf
        test_values[1] = 1.0; test_values[2] = 2.0; test_values[3] = 3.0;
        test_values[4] = 4.0; test_values[5] = 5.0; test_values[6] = 6.0; test_values[7] = 7.0;
        apply_test_case(test_values, neg_inf, "Test T16:  -Inf propagation", pass_count, fail_count);

        // 测试用例 17: Inf + (-Inf) = NaN
        test_values[0] = pos_inf; // +Inf
        test_values[1] = neg_inf; // -Inf
        test_values[2] = 1.0; test_values[3] = 2.0;
        test_values[4] = 3.0; test_values[5] = 4.0; test_values[6] = 5.0; test_values[7] = 6.0;
        apply_test_case(test_values, nan_val, "Test T17:  Inf + (-Inf) = NaN", pass_count, fail_count);

        // 测试用例 18: Inf + Inf = Inf
        test_values[0] = pos_inf; // +Inf
        test_values[1] = pos_inf; // +Inf
        test_values[2] = 1.0; test_values[3] = 2.0;
        test_values[4] = 3.0; test_values[5] = 4.0; test_values[6] = 5.0; test_values[7] = 6.0;
        apply_test_case(test_values, pos_inf, "Test T18:  Inf + Inf = Inf", pass_count, fail_count);

        // 测试用例 19: -Inf + -Inf = -Inf
        test_values[0] = neg_inf; // -Inf
        test_values[1] = neg_inf; // -Inf
        test_values[2] = 1.0; test_values[3] = 2.0;
        test_values[4] = 3.0; test_values[5] = 4.0; test_values[6] = 5.0; test_values[7] = 6.0;
        apply_test_case(test_values, neg_inf, "Test T19:  -Inf + -Inf = -Inf", pass_count, fail_count);

        // 测试用例 20: 多个 Inf (+/-) 混合 -> NaN
        test_values[0] = pos_inf; // +Inf
        test_values[1] = neg_inf; // -Inf
        test_values[2] = pos_inf; // +Inf
        test_values[3] = neg_inf; // -Inf
        test_values[4] = 1.0; test_values[5] = -1.0; test_values[6] = 0.0; test_values[7] = 0.0;
        apply_test_case(test_values, nan_val, "Test T20:  Multiple Inf (+/-) mix -> NaN", pass_count, fail_count);

        // 测试用例 21: 混合正零和负零 (预期结果为 +0.0)
        test_values[0] = 0.0; test_values[1] = -0.0; test_values[2] = 0.0; test_values[3] = -0.0;
        test_values[4] = 0.0; test_values[5] = -0.0; test_values[6] = 0.0; test_values[7] = -0.0;
        apply_test_case(test_values, 0.0, "Test T21:  Mixed +0 and -0 (expect +0)", pass_count, fail_count);

        // 测试用例 T22: 8个正零相加 (0 + 0 + ... + 0 = 0)
        test_values = '{0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0};
        apply_test_case(test_values, 0.0, "Table Test T22: 8 x +0", pass_count, fail_count);

        // 测试用例 T23: 8个负非规格化数相加
        test_values = '{-min_subnormal, -min_subnormal, -min_subnormal, -min_subnormal, -min_subnormal, -min_subnormal, -min_subnormal, -min_subnormal};
        expected_result = 8.0 * (-min_subnormal); // 结果为 -0.0 ：0x80000000见文档
        apply_test_case(test_values, expected_result, "Table Test T23: 8 x -denorm", pass_count, fail_count);

        // 测试用例 T24: 4个正非规格化数 + 4个负非规格化数 (相互抵消 = +0)
        test_values = '{min_subnormal, min_subnormal, min_subnormal, min_subnormal, -min_subnormal, -min_subnormal, -min_subnormal, -min_subnormal};
        apply_test_case(test_values, 0.0, "Table Test T24: 4 x +denorm + 4 x -denorm (Expect +0)", pass_count, fail_count);

        // 测试用例 T25: 8个 0x00800000 (最小正规格化数) 相加 
        // 8 * Val_00800000 = 8 * 2^-126 = 2^-123 (规格化数)
        test_values = '{val_00800000, val_00800000, val_00800000, val_00800000, val_00800000, val_00800000, val_00800000, val_00800000};
        expected_result = 8.0 * val_00800000;
        apply_test_case(test_values, expected_result, "Table Test T25: 8 x 0x00800000", pass_count, fail_count);

        // 测试用例 T26: 4个 +inf + 4个有限数
        test_values = '{pos_inf, pos_inf, pos_inf, pos_inf, 1.0, 2.0, 3.0, 4.0};
        apply_test_case(test_values, pos_inf, "Table Test T26: 4 x +inf + 4 x finite", pass_count, fail_count);

        // 测试用例 T27: 4个 -inf + 4个有限数
        test_values = '{neg_inf, neg_inf, neg_inf, neg_inf, 1.0, 2.0, 3.0, 4.0};
        apply_test_case(test_values, neg_inf, "Table Test T27: 4 x -inf + 4 x finite", pass_count, fail_count);

        // 测试用例 T28: 4个 +inf + 4个 -inf (结果为 NaN)
        test_values = '{pos_inf, pos_inf, pos_inf, pos_inf, neg_inf, neg_inf, neg_inf, neg_inf};
        apply_test_case(test_values, nan_val, "Table Test T28: 4 x +inf + 4 x -inf (Expect NaN)", pass_count, fail_count);

        // 测试用例 T29: 1个 NaN + 7个有限数 (结果为 NaN)
        test_values = '{nan_val, 1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0};
        apply_test_case(test_values, nan_val, "Table Test T29: 1 x NaN + 7 x finite (Expect NaN)", pass_count, fail_count);

        // 测试用例 T30: 1个 NaN + 7个 Inf (结果为 NaN)
        test_values = '{nan_val, pos_inf, neg_inf, pos_inf, neg_inf, pos_inf, neg_inf, pos_inf};
        apply_test_case(test_values, nan_val, "Table Test T30: 1 x NaN + 7 x Inf (Expect NaN)", pass_count, fail_count);

        // 测试用例 T31: 混合 Inf, NaN, 有限数 (结果为 NaN)
        test_values = '{pos_inf, neg_inf, nan_val, 1.0, -2.0, 0.0, min_subnormal, val_00800000};
        apply_test_case(test_values, nan_val, "Table Test T31: Mixed Inf, NaN, finite (Expect NaN)", pass_count, fail_count);

        // 测试用例 T32: 4个 0x007fffff + 4个 0x00800000 相加
        test_values = '{val_007fffff, val_007fffff, val_007fffff, val_007fffff, val_00800000, val_00800000, val_00800000, val_00800000};
        expected_result = 4.0 * val_00800000;
        apply_test_case(test_values, expected_result, "Table Test T32: 4 x 0x007fffff + 4 x 0x00800000", pass_count, fail_count);

        // 测试用例 T33: 0x007fffff + 0x00800000 (pairwise from table, extended to 8 inputs with zeros)
        test_values = '{val_007fffff, val_00800000, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0};
        expected_result = val_00800000;
        apply_test_case(test_values, expected_result, "Table Test T33: 0x007fffff + 0x00800000 (pairwise test)", pass_count, fail_count);

        // 测试用例 T34: 8 x 1.23
        test_values = '{1.23, 1.23, 1.23, 1.23, 1.23, 1.23, 1.23, 1.23};
        expected_result = 8.0 * 1.23;
        apply_test_case(test_values, expected_result, "Arbitrary Test T34: 8 x 1.23", pass_count, fail_count);

        // 测试用例 T35: 8 x -4.56
        test_values = '{-4.56, -4.56, -4.56, -4.56, -4.56, -4.56, -4.56, -4.56};
        expected_result = 8.0 * (-4.56);
        apply_test_case(test_values, expected_result, "Arbitrary Test T35: 8 x -4.56", pass_count, fail_count);

        // 测试用例 T36: 小量级正数相加 (1e-5 + 2e-5 + ... + 8e-5)
        test_values = '{1e-5, 2e-5, 3e-5, 4e-5, 5e-5, 6e-5, 7e-5, 8e-5};
        expected_result = (1.0+2.0+3.0+4.0+5.0+6.0+7.0+8.0) * 1e-5; // 结果为 3.6e-4
        apply_test_case(test_values, expected_result, "Arbitrary Test T36: Sum of small positive numbers", pass_count, fail_count);

        // 测试用例 T37: 大量级正数相加 (1e5 + 2e5 + ... + 8e5)
        test_values = '{1e5, 2e5, 3e5, 4e5, 5e5, 6e5, 7e5, 8e5};
        expected_result = (1.0+2.0+3.0+4.0+5.0+6.0+7.0+8.0) * 1e5; // 结果为 3.6e6
        apply_test_case(test_values, expected_result, "Arbitrary Test T37: Sum of large positive numbers", pass_count, fail_count);

        // 测试用例 T38: 混合量级和符号的数相加
        test_values = '{1.234, 5.678e-2, -9.012e3, 3.456, -1.234, -5.678e-2, 9.012e3, -3.456};
        expected_result = 0.0 ;// 结果为 0.0
        apply_test_case(test_values, expected_result, "Arbitrary Test T38: Mixed magnitude and sign numbers", pass_count, fail_count);

        // 测试用例 T39: 精确小数相加 (0.125 + 0.25 + ...)
        test_values = '{0.125, 0.25, 0.375, 0.5, 0.625, 0.75, 0.875, 1.0};
        expected_result = 0.125 + 0.25 + 0.375 + 0.5 + 0.625 + 0.75 + 0.875 + 1.0; // 结果为 4.5
        apply_test_case(test_values, expected_result, "Arbitrary Test T39: Sum of precise decimals", pass_count, fail_count);

        // 测试用例 T40: 正负数相加 (1.1 + -2.2 + 3.3 + -4.4 + 5.5 + -6.6 + 7.7 + -8.8)
        test_values = '{1.1, -2.2, 3.3, -4.4, 5.5, -6.6, 7.7, -8.8};
        expected_result = 1.1 + -2.2 + 3.3 + -4.4 + 5.5 + -6.6 + 7.7 + -8.8; // 结果为 -4.4
        apply_test_case(test_values, expected_result, "Arbitrary Test T40: Mixed positive and negative numbers", pass_count, fail_count);

        /*
        ***直接输入二进制数
        **/
        // 测试用例 T41: 8个 0x80000000 (-0.0) 相加
        for (int k=0; k<NUM_INPUTS; k++) hex_input_values_neg_zero[k] = 32'h80000000;
        expected_hex_sum_pos_zero = 32'h80000000; // 期望 -0.0 (0x80000000)
        apply_test_case_hex_inputs(hex_input_values_neg_zero, expected_hex_sum_pos_zero, "Test T41:  Direct Hex: 8 x -0.0 (0x80000000) ", pass_count, fail_count);

        // 测试用例 T42: 8 个最小正非规格化数 (0x00000001)
        for (int k = 0; k < NUM_INPUTS; k++) hex_inputs_min_subnormal[k] = 32'h00000001;
        expected_sum_min_subnormal = 32'h00000008; // 8 * 0x00000001 = 0x00000008
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T42: Direct Hex: 8 x 0x00000001", pass_count, fail_count);
        // 测试用例 T43: 8 个最大正非规格化数 (0x007FFFFF)
        for (int k = 0; k < NUM_INPUTS; k++) hex_inputs_max_subnormal[k] = 32'h007FFFFF;
        expected_sum_max_subnormal = 32'h01fFFFFE; // 已校正的最大非规格化数之和
        apply_test_case_hex_inputs(hex_inputs_max_subnormal, expected_sum_max_subnormal, "Test T43: Direct Hex: 8 x 0x007FFFFF", pass_count, fail_count);
        // 测试用例 T44: 8 个两倍最小正非规格化数 (0x00000002)
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            hex_inputs_min_subnormal[i] = 32'h00000002; // 8 * (2 * 2^-149)
        end
        expected_sum_min_subnormal = 32'h00000010; // 16 * 2^-149
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T44: Direct Hex: 8 x 0x00000002", pass_count, fail_count);

        // Test T45: 8 x 0x00000001 (smallest positive denormalized)
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            hex_inputs_min_subnormal[i] = 32'h00000001; // 8 * (1 * 2^-149)
        end
        expected_sum_min_subnormal = 32'h00000008;    // 8 * 2^-149
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T45: Direct Hex: 8 x 0x00000001", pass_count, fail_count);

        // Test T46: 4 x 0x00000001 + 4 x 0x00000002
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            if (i < 4) hex_inputs_min_subnormal[i] = 32'h00000001; // 4 * (1 * 2^-149)
            else       hex_inputs_min_subnormal[i] = 32'h00000002; // 4 * (2 * 2^-149)
        end
        expected_sum_min_subnormal = 32'h0000000C;
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T46: Direct Hex: 4x0x00000001 + 4x0x00000002", pass_count, fail_count);

        // Test T47: 2 x 0x00000003 + 2 x 0x00000004 + 4 x 0x00000001
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            if (i < 2)       hex_inputs_min_subnormal[i] = 32'h00001003; // 2 * (3 * 2^-149)
            else if (i < 4)  hex_inputs_min_subnormal[i] = 32'h00003004; // 2 * (4 * 2^-149)
            else             hex_inputs_min_subnormal[i] = 32'h0000f001; // 4 * (1 * 2^-149)
        end
        expected_sum_min_subnormal = 32'h00044012;
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T47: Direct Hex: 2x0x03 + 2x0x04 + 4x0x01", pass_count, fail_count);

        // Test T48: Sum resulting in a larger denormalized number (e.g., 8 x 0x00000010)
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            hex_inputs_min_subnormal[i] = 32'h00000010; // 8 * (16 * 2^-149)
        end
        expected_sum_min_subnormal = 32'h00000080;
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T48: Direct Hex: 8 x 0x00000010", pass_count, fail_count);

        // Test T49: Sum of denormalized numbers that could potentially normalize (e.g., 8 x 0x00100000)
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            hex_inputs_min_subnormal[i] = 32'h00100000;
        end
        expected_sum_min_subnormal = 32'h00800000; // Smallest positive normal number
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T49: Denorm sum to smallest Normal: 8 x 0x00100000", pass_count, fail_count);
        
        // Test T50: 8 x 0x00100001 (denormalized) resulting in a normal number
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            hex_inputs_min_subnormal[i] = 32'h00100001;
        end
        expected_sum_min_subnormal = 32'h00800008; // (1.00000000000000000000100)_2 * 2^-126
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T50: Denorm sum to Normal: 8 x 0x00100001", pass_count, fail_count);

        // Test T51: Alternating small denormalized numbers 0x00000001 and 0x00000002
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            if (i % 2 == 0) hex_inputs_min_subnormal[i] = 32'h00000001;
            else            hex_inputs_min_subnormal[i] = 32'h00000002;
        end
        expected_sum_min_subnormal = 32'h0000000C;
        apply_test_case_hex_inputs(hex_inputs_min_subnormal, expected_sum_min_subnormal, "Test T51: Alternating 0x01 and 0x02", pass_count, fail_count);
        
        // Test T52: 8 x Max Denormalized (0x007FFFFF)
        for (i = 0; i < NUM_INPUTS; i = i + 1) begin
            hex_inputs_max_subnormal[i] = 32'h007FFFFF;
        end
        expected_sum_max_subnormal = 32'h01FFFFFE; 
        apply_test_case_hex_inputs(hex_inputs_max_subnormal, 32'h01FFFFFE, "Test T52: 8 x Max Denormalized (0x007FFFFF)", pass_count, fail_count);

        // --- End of Additional Denormalized Number Test Cases ---



    // 显示测试结果统计
        $display("\n--- Test Summary ---");
        $display("Total PASS: %0d", pass_count);
        $display("Total FAIL: %0d", fail_count);
        
        $fdisplay(log_file, "\n--- Test Summary ---");
        $fdisplay(log_file, "Total PASS: %0d", pass_count);
        $fdisplay(log_file, "Total FAIL: %0d", fail_count);
        
        // 关闭日志文件
        $fclose(log_file);
        #(CLK_PERIOD * 10);
        $finish; // 结束仿真
    end


endmodule
